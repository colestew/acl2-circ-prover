<circuit>
    <CurrentPage>0</CurrentPage>
    <page 0>
    <PageViewport>-80.8805,16.9148,85.2529,-82.1518</PageViewport>
    <gate>
        <ID>16</ID>
        <type>AA_AND3</type>
        <position>-22.5,-7.5</position>
        <input>
            <ID>IN_0</ID>22
        </input>
        <input>
            <ID>IN_1</ID>18
        </input>
        <input>
            <ID>IN_2</ID>20
        </input>
        <output>
            <ID>OUT</ID>1
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 3</lparam>
    </gate>
    <gate>
        <ID>18</ID>
        <type>AA_AND3</type>
        <position>-23.5,-18</position>
        <input>
            <ID>IN_0</ID>20
        </input>
        <input>
            <ID>IN_1</ID>21
        </input>
        <input>
            <ID>IN_2</ID>19
        </input>
        <output>
            <ID>OUT</ID>2
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 3</lparam>
    </gate>
    <gate>
        <ID>26</ID>
        <type>BE_NOR3</type>
        <position>-4.5,-38.5</position>
        <input>
            <ID>IN_0</ID>6
        </input>
        <input>
            <ID>IN_1</ID>7
        </input>
        <input>
            <ID>IN_2</ID>20
        </input>
        <output>
            <ID>OUT</ID>5
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 3</lparam>
    </gate>
    <gate>
        <ID>28</ID>
        <type>BE_NOR2</type>
        <position>-7,-13.5</position>
        <input>
            <ID>IN_0</ID>1
        </input>
        <input>
            <ID>IN_1</ID>2
        </input>
        <output>
            <ID>OUT</ID>8
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 2</lparam>
    </gate>
    <gate>
        <ID>30</ID>
        <type>AA_AND2</type>
        <position>15.5,-2.5</position>
        <input>
            <ID>IN_0</ID>8
        </input>
        <output>
            <ID>OUT</ID>10
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 2</lparam>
    </gate>
    <gate>
        <ID>32</ID>
        <type>AA_AND3</type>
        <position>16,-9.5</position>
        <input>
            <ID>IN_0</ID>8
        </input>
        <output>
            <ID>OUT</ID>11
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 3</lparam>
    </gate>
    <gate>
        <ID>34</ID>
        <type>BE_NOR4</type>
        <position>33.5,-9</position>
        <input>
            <ID>IN_0</ID>5
        </input>
        <input>
            <ID>IN_1</ID>10
        </input>
        <input>
            <ID>IN_2</ID>11
        </input>
        <input>
            <ID>IN_3</ID>12
        </input>
        <output>
            <ID>OUT</ID>9
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 4</lparam>
    </gate>
    <gate>
        <ID>36</ID>
        <type>AA_AND4</type>
        <position>16,-17</position>
        <input>
            <ID>IN_0</ID>8
        </input>
        <output>
            <ID>OUT</ID>12
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 4</lparam>
    </gate>
    <gate>
        <ID>44</ID>
        <type>AA_AND2</type>
        <position>-23.5,-35</position>
        <input>
            <ID>IN_0</ID>19
        </input>
        <input>
            <ID>IN_1</ID>26
        </input>
        <output>
            <ID>OUT</ID>6
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 2</lparam>
    </gate>
    <gate>
        <ID>46</ID>
        <type>AA_AND2</type>
        <position>-23.5,-42</position>
        <input>
            <ID>IN_0</ID>27
        </input>
        <input>
            <ID>IN_1</ID>22
        </input>
        <output>
            <ID>OUT</ID>7
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 2</lparam>
    </gate>
    <gate>
        <ID>48</ID>
        <type>AI_XOR2</type>
        <position>17.5,-48</position>
        <input>
            <ID>IN_0</ID>8
        </input>
        <input>
            <ID>IN_1</ID>5
        </input>
        <output>
            <ID>OUT</ID>4
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 2</lparam>
    </gate>
    <gate>
        <ID>50</ID>
        <type>DI_NAND8</type>
        <position>16,-26</position>
        <input>
            <ID>IN_0</ID>8
        </input>
        <output>
            <ID>OUT</ID>13
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 8</lparam>
    </gate>
    <gate>
        <ID>52</ID>
        <type>BA_NAND4</type>
        <position>16.5,-35</position>
        <input>
            <ID>IN_0</ID>8
        </input>
        <output>
            <ID>OUT</ID>23
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 4</lparam>
    </gate>
    <gate>
        <ID>54</ID>
        <type>AI_XOR2</type>
        <position>47.5,-49</position>
        <input>
            <ID>IN_0</ID>4
        </input>
        <output>
            <ID>OUT</ID>25
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 2</lparam>
    </gate>
    <gate>
        <ID>56</ID>
        <type>BI_NANDX2</type>
        <position>55,-23.5</position>
        <input>
            <ID>IN_0</ID>9
        </input>
        <input>
            <ID>IN_1</ID>13
        </input>
        <output>
            <ID>OUT</ID>24
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 2</lparam>
    </gate>
    <gate>
        <ID>68</ID>
        <type>DA_FROM</type>
        <position>-66,8</position>
        <input>
            <ID>IN_0</ID>18
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID S3</lparam>
    </gate>
    <gate>
        <ID>70</ID>
        <type>DA_FROM</type>
        <position>-66,4.5</position>
        <input>
            <ID>IN_0</ID>21
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID S2</lparam>
    </gate>
    <gate>
        <ID>72</ID>
        <type>DA_FROM</type>
        <position>-66.5,0.5</position>
        <input>
            <ID>IN_0</ID>26
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID S1</lparam>
    </gate>
    <gate>
        <ID>74</ID>
        <type>DA_FROM</type>
        <position>-66.5,-3</position>
        <input>
            <ID>IN_0</ID>27
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID S0</lparam>
    </gate>
    <gate>
        <ID>76</ID>
        <type>DA_FROM</type>
        <position>-76,-24.5</position>
        <input>
            <ID>IN_0</ID>22
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID B3</lparam>
    </gate>
    <gate>
        <ID>78</ID>
        <type>DA_FROM</type>
        <position>-75.5,-48</position>
        <input>
            <ID>IN_0</ID>20
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID A3</lparam>
    </gate>
    <gate>
        <ID>82</ID>
        <type>AA_INVERTER</type>
        <position>-62.5,-24.5</position>
        <input>
            <ID>IN_0</ID>22
        </input>
        <output>
            <ID>OUT_0</ID>19
        </output>
        <gparam>angle 0.0</gparam>
        <lparam>INPUT_BITS 1</lparam>
    </gate>
    <gate>
        <ID>84</ID>
        <type>DE_TO</type>
        <position>73.5,-9</position>
        <input>
            <ID>IN_0</ID>9
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID Y</lparam>
    </gate>
    <gate>
        <ID>88</ID>
        <type>DE_TO</type>
        <position>75,-34.5</position>
        <input>
            <ID>IN_0</ID>23
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID X</lparam>
    </gate>
    <gate>
        <ID>90</ID>
        <type>DE_TO</type>
        <position>73.5,-48.5</position>
        <input>
            <ID>IN_0</ID>25
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID F3</lparam>
    </gate>
    <gate>
        <ID>92</ID>
        <type>DE_TO</type>
        <position>73.5,-24.5</position>
        <input>
            <ID>IN_0</ID>24
        </input>
        <gparam>angle 0.0</gparam>
        <lparam>JUNCTION_ID Cnot_p4</lparam>
    </gate>
    <wire>
        <ID>1</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-15,-12.5,-15,-7.5</points>
                <intersection>-12.5 1</intersection>
                <intersection>-7.5 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-15,-12.5,-10,-12.5</points>
                <connection>
                    <GID>28</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-15 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-19.5,-7.5,-15,-7.5</points>
                <connection>
                    <GID>16</GID>
                    <name>OUT</name>
                </connection>
                <intersection>-15 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>2</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-15,-18,-15,-14.5</points>
                <intersection>-18 2</intersection>
                <intersection>-14.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-15,-14.5,-10,-14.5</points>
                <connection>
                    <GID>28</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>-15 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-20.5,-18,-15,-18</points>
                <connection>
                    <GID>18</GID>
                    <name>OUT</name>
                </connection>
                <intersection>-15 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>4</ID>
        <shape>
            <hsegment>
                <ID>1</ID>
                <points>20.5,-48,44.5,-48</points>
                <connection>
                    <GID>48</GID>
                    <name>OUT</name>
                </connection>
                <connection>
                    <GID>54</GID>
                    <name>IN_0</name>
                </connection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>5</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-0.5,-49,-0.5,1.5</points>
                <intersection>-49 4</intersection>
                <intersection>-38.5 2</intersection>
                <intersection>1.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-0.5,1.5,30.5,1.5</points>
                <intersection>-0.5 0</intersection>
                <intersection>30.5 3</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-1.5,-38.5,-0.5,-38.5</points>
                <connection>
                    <GID>26</GID>
                    <name>OUT</name>
                </connection>
                <intersection>-0.5 0</intersection>
            </hsegment>
            <vsegment>
                <ID>3</ID>
                <points>30.5,-6,30.5,1.5</points>
                <connection>
                    <GID>34</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>1.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>4</ID>
                <points>-0.5,-49,14.5,-49</points>
                <connection>
                    <GID>48</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>-0.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>6</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-14,-36.5,-14,-35</points>
                <intersection>-36.5 1</intersection>
                <intersection>-35 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-14,-36.5,-7.5,-36.5</points>
                <connection>
                    <GID>26</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-14 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-20.5,-35,-14,-35</points>
                <connection>
                    <GID>44</GID>
                    <name>OUT</name>
                </connection>
                <intersection>-14 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>7</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-14,-42,-14,-38.5</points>
                <intersection>-42 2</intersection>
                <intersection>-38.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-14,-38.5,-7.5,-38.5</points>
                <connection>
                    <GID>26</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>-14 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-20.5,-42,-14,-42</points>
                <connection>
                    <GID>46</GID>
                    <name>OUT</name>
                </connection>
                <intersection>-14 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>8</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>5,-47,5,-1.5</points>
                <intersection>-47 1</intersection>
                <intersection>-32 8</intersection>
                <intersection>-22.5 7</intersection>
                <intersection>-14 4</intersection>
                <intersection>-13.5 2</intersection>
                <intersection>-1.5 3</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>5,-47,14.5,-47</points>
                <connection>
                    <GID>48</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-4,-13.5,5,-13.5</points>
                <connection>
                    <GID>28</GID>
                    <name>OUT</name>
                </connection>
                <intersection>5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>3</ID>
                <points>5,-1.5,12.5,-1.5</points>
                <connection>
                    <GID>30</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>5 0</intersection>
                <intersection>7 5</intersection>
            </hsegment>
            <hsegment>
                <ID>4</ID>
                <points>5,-14,13,-14</points>
                <connection>
                    <GID>36</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>5 0</intersection>
            </hsegment>
            <vsegment>
                <ID>5</ID>
                <points>7,-7.5,7,-1.5</points>
                <intersection>-7.5 6</intersection>
                <intersection>-1.5 3</intersection>
            </vsegment>
            <hsegment>
                <ID>6</ID>
                <points>7,-7.5,13,-7.5</points>
                <connection>
                    <GID>32</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>7 5</intersection>
            </hsegment>
            <hsegment>
                <ID>7</ID>
                <points>5,-22.5,13,-22.5</points>
                <connection>
                    <GID>50</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>8</ID>
                <points>5,-32,13.5,-32</points>
                <connection>
                    <GID>52</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>9</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>44.5,-9.5,44.5,-9</points>
                <intersection>-9.5 1</intersection>
                <intersection>-9 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>44.5,-9.5,71.5,-9.5</points>
                <intersection>44.5 0</intersection>
                <intersection>48 6</intersection>
                <intersection>71.5 5</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>37.5,-9,44.5,-9</points>
                <connection>
                    <GID>34</GID>
                    <name>OUT</name>
                </connection>
                <intersection>44.5 0</intersection>
            </hsegment>
            <vsegment>
                <ID>5</ID>
                <points>71.5,-9.5,71.5,-9</points>
                <connection>
                    <GID>84</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-9.5 1</intersection>
            </vsegment>
            <vsegment>
                <ID>6</ID>
                <points>48,-22.5,48,-9.5</points>
                <intersection>-22.5 7</intersection>
                <intersection>-9.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>7</ID>
                <points>48,-22.5,52,-22.5</points>
                <connection>
                    <GID>56</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>48 6</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>10</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>24.5,-8,24.5,-2.5</points>
                <intersection>-8 1</intersection>
                <intersection>-2.5 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>24.5,-8,30.5,-8</points>
                <connection>
                    <GID>34</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>24.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>18.5,-2.5,24.5,-2.5</points>
                <connection>
                    <GID>30</GID>
                    <name>OUT</name>
                </connection>
                <intersection>24.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>11</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>24.5,-10,24.5,-9.5</points>
                <intersection>-10 1</intersection>
                <intersection>-9.5 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>24.5,-10,30.5,-10</points>
                <connection>
                    <GID>34</GID>
                    <name>IN_2</name>
                </connection>
                <intersection>24.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>19,-9.5,24.5,-9.5</points>
                <connection>
                    <GID>32</GID>
                    <name>OUT</name>
                </connection>
                <intersection>24.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>12</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>24.5,-17,24.5,-12</points>
                <intersection>-17 2</intersection>
                <intersection>-12 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>24.5,-12,30.5,-12</points>
                <connection>
                    <GID>34</GID>
                    <name>IN_3</name>
                </connection>
                <intersection>24.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>19,-17,24.5,-17</points>
                <connection>
                    <GID>36</GID>
                    <name>OUT</name>
                </connection>
                <intersection>24.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>13</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>35.5,-26,35.5,-24.5</points>
                <intersection>-26 2</intersection>
                <intersection>-24.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>35.5,-24.5,52,-24.5</points>
                <connection>
                    <GID>56</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>35.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>19,-26,35.5,-26</points>
                <connection>
                    <GID>50</GID>
                    <name>OUT</name>
                </connection>
                <intersection>35.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>18</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-45,-7.5,-45,8</points>
                <intersection>-7.5 2</intersection>
                <intersection>8 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-64,8,-45,8</points>
                <connection>
                    <GID>68</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-45 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-45,-7.5,-25.5,-7.5</points>
                <connection>
                    <GID>16</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>-45 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>19</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-28.5,-34,-28.5,-20</points>
                <intersection>-34 4</intersection>
                <intersection>-24.5 1</intersection>
                <intersection>-20 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-59.5,-24.5,-28.5,-24.5</points>
                <connection>
                    <GID>82</GID>
                    <name>OUT_0</name>
                </connection>
                <intersection>-28.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-28.5,-20,-26.5,-20</points>
                <connection>
                    <GID>18</GID>
                    <name>IN_2</name>
                </connection>
                <intersection>-28.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>4</ID>
                <points>-28.5,-34,-26.5,-34</points>
                <connection>
                    <GID>44</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-28.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>20</ID>
        <shape>
            <hsegment>
                <ID>1</ID>
                <points>-73.5,-48.5,-7.5,-48.5</points>
                <intersection>-73.5 6</intersection>
                <intersection>-40 3</intersection>
                <intersection>-7.5 8</intersection>
            </hsegment>
            <vsegment>
                <ID>3</ID>
                <points>-40,-48.5,-40,-9.5</points>
                <intersection>-48.5 1</intersection>
                <intersection>-16 10</intersection>
                <intersection>-9.5 7</intersection>
            </vsegment>
            <vsegment>
                <ID>6</ID>
                <points>-73.5,-48.5,-73.5,-48</points>
                <connection>
                    <GID>78</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-48.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>7</ID>
                <points>-40,-9.5,-25.5,-9.5</points>
                <connection>
                    <GID>16</GID>
                    <name>IN_2</name>
                </connection>
                <intersection>-40 3</intersection>
            </hsegment>
            <vsegment>
                <ID>8</ID>
                <points>-7.5,-48.5,-7.5,-40.5</points>
                <connection>
                    <GID>26</GID>
                    <name>IN_2</name>
                </connection>
                <intersection>-48.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>10</ID>
                <points>-40,-16,-26.5,-16</points>
                <connection>
                    <GID>18</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-40 3</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>21</ID>
        <shape>
            <hsegment>
                <ID>1</ID>
                <points>-47,-18,-26.5,-18</points>
                <connection>
                    <GID>18</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>-47 3</intersection>
            </hsegment>
            <vsegment>
                <ID>3</ID>
                <points>-47,-18,-47,4.5</points>
                <intersection>-18 1</intersection>
                <intersection>4.5 4</intersection>
            </vsegment>
            <hsegment>
                <ID>4</ID>
                <points>-64,4.5,-47,4.5</points>
                <connection>
                    <GID>70</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-47 3</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>22</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-71,-43,-71,-5.5</points>
                <intersection>-43 4</intersection>
                <intersection>-24.5 1</intersection>
                <intersection>-24.5 1</intersection>
                <intersection>-5.5 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-74,-24.5,-65.5,-24.5</points>
                <connection>
                    <GID>76</GID>
                    <name>IN_0</name>
                </connection>
                <connection>
                    <GID>82</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-71 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-71,-5.5,-25.5,-5.5</points>
                <connection>
                    <GID>16</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-71 0</intersection>
            </hsegment>
            <hsegment>
                <ID>4</ID>
                <points>-71,-43,-26.5,-43</points>
                <connection>
                    <GID>46</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>-71 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>23</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>46,-35,46,-34.5</points>
                <intersection>-35 2</intersection>
                <intersection>-34.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>46,-34.5,73,-34.5</points>
                <connection>
                    <GID>88</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>46 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>19.5,-35,46,-35</points>
                <connection>
                    <GID>52</GID>
                    <name>OUT</name>
                </connection>
                <intersection>46 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>24</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>64.5,-24.5,64.5,-23.5</points>
                <intersection>-24.5 1</intersection>
                <intersection>-23.5 2</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>64.5,-24.5,71.5,-24.5</points>
                <connection>
                    <GID>92</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>64.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>58,-23.5,64.5,-23.5</points>
                <connection>
                    <GID>56</GID>
                    <name>OUT</name>
                </connection>
                <intersection>64.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>25</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>61,-49,61,-48.5</points>
                <intersection>-49 2</intersection>
                <intersection>-48.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>61,-48.5,71.5,-48.5</points>
                <connection>
                    <GID>90</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>61 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>50.5,-49,61,-49</points>
                <connection>
                    <GID>54</GID>
                    <name>OUT</name>
                </connection>
                <intersection>61 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>26</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-49,-36,-49,0.5</points>
                <intersection>-36 2</intersection>
                <intersection>0.5 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-64.5,0.5,-49,0.5</points>
                <connection>
                    <GID>72</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-49 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-49,-36,-26.5,-36</points>
                <connection>
                    <GID>44</GID>
                    <name>IN_1</name>
                </connection>
                <intersection>-49 0</intersection>
            </hsegment>
        </shape>
    </wire>
    <wire>
        <ID>27</ID>
        <shape>
            <vsegment>
                <ID>0</ID>
                <points>-51.5,-41,-51.5,-3</points>
                <intersection>-41 2</intersection>
                <intersection>-3 1</intersection>
            </vsegment>
            <hsegment>
                <ID>1</ID>
                <points>-64.5,-3,-51.5,-3</points>
                <connection>
                    <GID>74</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-51.5 0</intersection>
            </hsegment>
            <hsegment>
                <ID>2</ID>
                <points>-51.5,-41,-26.5,-41</points>
                <connection>
                    <GID>46</GID>
                    <name>IN_0</name>
                </connection>
                <intersection>-51.5 0</intersection>
            </hsegment>
        </shape>
    </wire>
    </page 0>
    <page 1>
    <PageViewport>-80.8805,16.9148,85.2529,-82.1518</PageViewport>
    </page 1>
    <page 2>
    <PageViewport>-80.8805,16.9148,85.2529,-82.1518</PageViewport>
    </page 2>
    <page 3>
    <PageViewport>-80.8805,16.9148,85.2529,-82.1518</PageViewport>
    </page 3>
    <page 4>
    <PageViewport>-80.8805,16.9148,85.2529,-82.1518</PageViewport>
    </page 4>
    <PageViewport>-80.8805,16.9148,85.2529,-82.1518</PageViewport>
    </page >

</circuit>
